-- Secondary GR1553B
  constant CFG_GR1553B_ENABLE2    : integer := CONFIG_GR1553B_ENABLE2;
  constant CFG_GR1553B_RTEN2      : integer := CONFIG_GR1553B_RTEN2;
  constant CFG_GR1553B_BCEN2      : integer := CONFIG_GR1553B_BCEN2;
  constant CFG_GR1553B_BMEN2      : integer := CONFIG_GR1553B_BMEN2;
