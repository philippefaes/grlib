
package DW_Foundation_arith is

end;
