-- PCIEXP	interface
	constant CFG_PCIEXP         : integer	:= CFG_PCIE;
	constant CFG_PCIE_TYPE			:	integer	:= CFG_PCIETYPE;
	constant CFG_PCIE_SIM_MAS		:	integer	:= CFG_PCIEMASTER;
	constant CFG_PCIEXPVID			:	integer	:= 16#CONFIG_PCIEXP_VENDORID#;
	constant CFG_PCIEXPDID			:	integer	:= 16#CONFIG_PCIEXP_DEVICEID#;
  constant CFG_NO_OF_LANES    : integer := CFG_LANE_WIDTH;
