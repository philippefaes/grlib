-- SPI to AHB bridge
  constant CFG_SPI2AHB         : integer := CONFIG_SPI2AHB;
  constant CFG_SPI2AHB_APB     : integer := CONFIG_SPI2AHB_APB;
  constant CFG_SPI2AHB_ADDRH   : integer := 16#CONFIG_SPI2AHB_ADDRH#;
  constant CFG_SPI2AHB_ADDRL   : integer := 16#CONFIG_SPI2AHB_ADDRL#;
  constant CFG_SPI2AHB_MASKH   : integer := 16#CONFIG_SPI2AHB_MASKH#;
  constant CFG_SPI2AHB_MASKL   : integer := 16#CONFIG_SPI2AHB_MASKL#;
  constant CFG_SPI2AHB_RESEN   : integer := CONFIG_SPI2AHB_RESEN;
  constant CFG_SPI2AHB_FILTER  : integer := CONFIG_SPI2AHB_FILTER;
  constant CFG_SPI2AHB_CPOL    : integer := CONFIG_SPI2AHB_CPOL;
  constant CFG_SPI2AHB_CPHA    : integer := CONFIG_SPI2AHB_CPHA;
